
/******************************************************************************/
// `include "gParam.v"
//==============================================================================
`timescale 1ns/100ps

`include "RTL/PLL.v"
//==============================================================================
module PLL_tb;
//------------------------------------------------------------------------------
//  UUT
//------------------------------------------------------------------------------
    // ports
    reg     RST     ;  // 
    reg     CLK     ;  // 
    wire    CLK45   ;  // 
    wire    CLK90   ;  // 
    wire    CLK135  ;  // 
    wire    LOCKED  ;  // 
    // module
    PLL uut (
        .RST        (RST      ),
        .CLK        (CLK      ),
        .CLK45      (CLK45    ),
        .CLK90      (CLK90    ),
        .CLK135     (CLK135   ),
        .LOCKED     (LOCKED   )
    );
//------------------------------------------------------------------------------
//  localparam
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
//  clk
//------------------------------------------------------------------------------
    localparam CLK_FREQ = 25_000_000;
    localparam PERIOD = 1E9/CLK_FREQ;
    initial begin
        CLK = 0;
        forever #(PERIOD/2) CLK = ~ CLK;
    end
//------------------------------------------------------------------------------
//  general tasks and functions
//------------------------------------------------------------------------------
    // -------- wait n periods of clock --------
    task wait_n_clk(input integer i);
        begin
            repeat(i) @(posedge CLK);
        end
    endtask
    // -------- wait n periods of clock (with Tcko) --------
    task wait_n_clko(input integer i);
        begin
            repeat(i) @(posedge CLK);
            #1;
        end
    endtask
//------------------------------------------------------------------------------
//  initial values
//------------------------------------------------------------------------------
    initial begin
        RST = 1;
        // -------- input --------
    end
//------------------------------------------------------------------------------
//  simulation tasks
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
//  run simulation
//------------------------------------------------------------------------------
    initial begin
        $display("*Testing PLL Mock for Simulation*");
        $dumpfile("../VCD/PLL_tb.vcd");
        $dumpvars(0, PLL_tb);
        // -------- RESET --------
        wait_n_clk(2);
        RST = 1;
        wait_n_clko(2);
        RST = 0;
        wait_n_clko(20);
        $finish;
    end
//------------------------------------------------------------------------------
endmodule