 /*
// 
// Copyright (C) 2022  Mike Taylor
// This file is part of RE-SDMAC <https://github.com/mbtaylor1982/RE-SDMAC>.
// 
// RE-SDMAC is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
// 
// RE-SDMAC is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with dogtag.  If not, see <http://www.gnu.org/licenses/>.
 */
module fifo_byte_ptr(
    input INCBO,
    input MID25,
    input ACR_WR,
    input H_0C,
    input RST_FIFO_,    

    output reg [1:0] PTR    
);

wire MUXZ;

always @(posedge ACR_WR or posedge INCBO or negedge RST_FIFO_) begin
    if (RST_FIFO_ == 1'b0) 
        PTR <= 2'b00;
    else begin
        if (INCBO) PTR <= {MUXZ, ~PTR[0]};
        if (ACR_WR) PTR[1] <= MUXZ;        
    end    
end

assign MUXZ = (H_0C)? ~MID25:(PTR[0]^~PTR[1]);

endmodule