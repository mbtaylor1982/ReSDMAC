
/******************************************************************************/
// `include "gParam.v"
//==============================================================================
`timescale 1ns/100ps

`include "RTL/PLL.v"
//==============================================================================
module PLL_tb;
//------------------------------------------------------------------------------
//  UUT
//------------------------------------------------------------------------------
    // ports
    reg     rst   ;  // 
    reg     CPUCLK_I   ;  // 
    wire    nCLK   ;  // 
    wire    BCLK   ;  // 
    wire    BBCLK  ;  // 
    wire    QnCPUCLK;
    wire    locked;  // 
    // module
    PLL uut (
        .RST        (rst      ),
        .CLK        (CPUCLK_I ),
        .CLK45      (nCLK     ),
        .CLK90      (BCLK     ),
        .CLK135     (BBCLK    ),
        .LOCKED     (locked   )
    );
//------------------------------------------------------------------------------
//  localparam
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
//  clk
//------------------------------------------------------------------------------
    localparam CLK_FREQ = 25_000_000;
    localparam PERIOD = 1E9/CLK_FREQ;
    initial begin
        CPUCLK_I = 0;
        forever #(PERIOD/2) CPUCLK_I = ~ CPUCLK_I;
    end
//------------------------------------------------------------------------------
//  general tasks and functions
//------------------------------------------------------------------------------
    // -------- wait n periods of clock --------
    task wait_n_clk(input integer i);
        begin
            repeat(i) @(posedge CPUCLK_I);
        end
    endtask
    // -------- wait n periods of clock (with Tcko) --------
    task wait_n_clko(input integer i);
        begin
            repeat(i) @(posedge CPUCLK_I);
            #1;
        end
    endtask
//------------------------------------------------------------------------------
//  initial values
//------------------------------------------------------------------------------
    initial begin
        rst = 1;
        // -------- input --------

    end
//------------------------------------------------------------------------------
//  simulation tasks
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
//  run simulation
//------------------------------------------------------------------------------
    initial begin
        $display("*Testing PLL Mock for Simulation*");
        $dumpfile("../VCD/PLL_tb.vcd");
        $dumpvars(0, PLL_tb);
        // -------- RESET --------
        wait_n_clk(2);
        rst = 1;
        wait_n_clko(2);
        rst = 0;
        wait_n_clko(20);
        $finish;
    end

    assign QnCPUCLK = ~CPUCLK_I;
//------------------------------------------------------------------------------
endmodule