/*
// 
// Copyright (C) 2022  Mike Taylor
// This file is part of RE-SDMAC <https://github.com/mbtaylor1982/RE-SDMAC>.
// 
// RE-SDMAC is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
// 
// RE-SDMAC is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with dogtag.  If not, see <http://www.gnu.org/licenses/>.
 */
module CPU_SM_outputs (
    input E32, E48,
    input E2, E3, E4, E5, E7, E8, 
    input E10, E11, E12, E16, E17, E18,
    input E19,
    input E0, E21, E26, E27,
    input E56, E55, E35, E61, E50_d_E52_d,
    input E60, DSACK, E43_s_E49_sd, E57_s, STERM_,
    input E36_s_E47_s, E33_sd_E38_s, E40_s_E41_s, E42_s, E46_s_E59_s, E51_s_E54_sd,
    input E62, E58, E53, E25_d, E28_d, E30_d,
    input E23_sd, E29_sd,
    input E45, E34, E24_sd, E37_s, E44_s,

    output nINCNI_d,
    output nBREQ_d,
    output SIZE1_d,
    output PAS_d,
    output PDS_d,
    output F2CPUL_d,
    output F2CPUH_d,
    output BRIDGEOUT_d,

    output PLLW_d,
    output PLHW_d,
    output INCFIFO_d,
    output DECFIFO_d,
    output INCNO_d,
    output nSTOPFLUSH_d,
    output DIEH_d,
    output DIEL_d,
    output nBRIDGEIN_d,
    output BGACK_d
);


assign nINCNI_d = (~(E32 | E48)); 
//assign INCNI_d = (E32 | E48);
assign nBREQ_d = (~((E2 | E3 | E4 | E5 | E7 | E8) | (E10 | E11 | E12 | E16 | E17 | E18) | E19)); 
//assign BREQ_d = ((E2 | E3 | E4 | E5 | E7 | E8) | (E10 | E11 | E12 | E16 | E17 | E18) | E19);


//SIZE1
wire SIZE1_X, SIZE1_Y, SIZE1_Z;

assign SIZE1_X = (~((~E62 & ~E61 & ~E58 & ~E56 & ~E53 & ~E26) & ~(~(~E25_d & ~E28_d & ~E30_d & ~E50_d_E52_d) & DSACK) & ~(E50_d_E52_d & ~DSACK)));
assign SIZE1_Y = (~(~STERM_ & ~(~E36_s_E47_s & ~E33_sd_E38_s & ~E40_s_E41_s & ~E42_s & ~E46_s_E59_s & ~E51_s_E54_sd)));
assign SIZE1_Z = (~((~(~(E23_sd & DSACK) & ~(~DSACK & (E29_sd | E33_sd_E38_s | E51_s_E54_sd))) |(E40_s_E41_s | E36_s_E47_s | E46_s_E59_s)) & STERM_));

assign SIZE1_d = (~(SIZE1_X & SIZE1_Y & SIZE1_Z));

//PAS
wire PAS_X, PAS_Y;
assign PAS_X = (~(~(~E62 & ~E61 & ~E60 & ~E58) |~(~E56 & ~E53 & ~E48 & ~E45) | ~(~E34 & ~E26 & ~E21)) & ~(E50_d_E52_d & ~DSACK));
assign PAS_Y = (~(((~DSACK & (E24_sd | E29_sd | E33_sd_E38_s | E43_s_E49_sd | E51_s_E54_sd))|(E37_s-E44_s | E40_s_E41_s | E36_s_E47_s | E57_s | E46_s_E59_s)) & STERM_));

assign PAS_d = (~(PAS_X & PAS_Y));

//assign PDS_d = ;
//assign F2CPUL_d = ; 
//assign F2CPUH_d = ;
//assign BRIDGEOUT_d = ;
//assign PLLW_d = ;
assign PLHW_d = ~(~(E48 | E60) & (~(((~DSACK & E43_s_E49_sd) | E57_s) & STERM_)));
//assign INCFIFO_d = ;
//assign DECFIFO_d = ;
//assign INCNO_d = ;
assign nSTOPFLUSH_d = (~E0 & ~E4 & ~E5 & ~E21 & ~E26 & ~E27); 
//assign STOPFLUSH_d = (E0 | E4 | E5 | E21 | E26 | E27);
//assign DIEH_d = ;
//assign DIEL_d = ;
assign nBRIDGEIN_d = (~(~E56 & ~E55 & ~E35 & ~E61 & ~E50_d_E52_d));
//assign BRIDGEIN_d = ~(E56 | E55 | E35 | E61 | E50_d_E52_d);
//assign BGACK_d = ;

endmodule